module top(
  input clk,
  input rst,
  input en_pb,
  output [3:0] vgaRed,
  output [3:0] vgaGreen,
  output [3:0] vgaBlue,
  output hsync,
  output vsync
);

wire [11:0] data;
wire clk_25MHz;
wire clk_22;
wire clk_100Hz;
wire [16:0] pixel_addr;
wire [11:0] pixel;
wire valid;
wire [9:0] h_cnt; //640
wire [9:0] v_cnt;  //480
wire en_debounced;
wire en_onepulse;
reg en_scroll,en_scroll_next;


assign {vgaRed, vgaGreen, vgaBlue} = (valid==1'b1) ? pixel:12'h0;


always@(posedge clk_22)
begin
    if(rst)
        en_scroll <= 1'b0;
     else
        en_scroll <= en_scroll_next;
end

always@*
begin
    en_scroll_next = 1'b0;
    case(en_scroll)
    1'b1: en_scroll_next = (en_onepulse == 1'b1)? 1'b0:1'b1;
    1'b0: en_scroll_next = (en_onepulse == 1'b1)? 1'b1:1'b0;
    endcase
end

// Frequency Divider
Frequency_Divider U0(
  .clk(clk),
  .rst_n(~rst), 
  .clk1(clk_25MHz),
  .clk_100Hz(clk_100Hz),
  .clk22(clk_22)
);


debounce_circuit U1(
    .clk(clk_100Hz), 
    .rst_n(~rst), 
    .pb_in(en_pb), 
    .pb_debounced(en_debounced)
);

one_pulse U2(
  .clk(clk_22), 
  .rst_n(~rst),
  .in_trig(en_pb), 
  .out_pulse(en_onepulse) 
);

// Reduce frame address from 640x480 to 320x240
mem_addr_gen mem_addr_gen_inst(
  .clk(clk_22),
  .rst(rst),
  .h_cnt(h_cnt),
  .v_cnt(v_cnt),
  .en_scroll(en_scroll),
  .pixel_addr(pixel_addr)
);
     
// Use reduced 320x240 address to output the saved picture from RAM 
blk_mem_gen_0 blk_mem_gen_0_inst(
  .clka(clk_25MHz),
  .wea(0),
  .addra(pixel_addr),
  .dina(data[11:0]),
  .douta(pixel)
); 

// Render the picture by VGA controller
vga_controller   vga_inst(
  .pclk(clk_25MHz),
  .reset(rst),
  .hsync(hsync),
  .vsync(vsync),
  .valid(valid),
  .h_cnt(h_cnt),
  .v_cnt(v_cnt)
);
      
endmodule
